module InstMem(addr, dout);
	input logic [4:0] addr;
	output logic [31:0] dout;
	bit [31:0] mem [35:0] = '{32'b00010000000000000000100100010111,
							  32'b0, 32'b0, 32'b0,
							  32'b00000000000010010000100100010011,
							  32'b0, 32'b0, 32'b0,
							  32'b00000000000010010010101000000011,
							  32'b0, 32'b0, 32'b0,
							  32'b00000000010010010010101010000011,
							  32'b0, 32'b0, 32'b0,
							  32'b00000001010110100000101000110011,
							  32'b0, 32'b0, 32'b0,
							  32'b01000001010110100000101010110011,
							  32'b0, 32'b0, 32'b0,
							  32'b01000001010110100000101000110011,
							  32'b0, 32'b0, 32'b0,
							  32'b00000001010010010010000000100011,
							  32'b0, 32'b0, 32'b0,
							  32'b00000001010110010010000000100011,
							  32'b0, 32'b0, 32'b0
							 };
	assign dout = mem[addr];
endmodule